------------------------------------
-- Class 3 Example 1: D/JK-FlipFlop
------------------------------------
-- Version: 1.0
-- Author: Max Gundacker
-- Date: 05 May 2025
-- Filename: FlipFlop_rtl_cfg.vhd
------------------------------------
-- Description: configuration of 
-- FlipFlop for example 1
------------------------------------

configuration counter_rtl_cfg of counter is
	for rtl
	end for;
end counter_rtl_cfg;
