-------------------------------------------------------------------
--          Microelectronic Design | FH Technikum Wien           --
--                        COUNTER PROJECT                        --
-------------------------------------------------------------------
--       Author: Bauer Julian  (el23b071@technikum-wien.at)      --
--               Gundacker Max (el23b074@technikum-wien.at)      --
--                                                               --
--         Date: 24 Jun 2025                                     --
--                                                               --
--  Design Unit: Counter Unit (Config)                           --
--                                                               --
--     Filename: counter_rtl_cfg.vhd                             --
--                                                               --
--      Version: 1.0                                             --
--                                                               --
--  Description: The counter unit implements a 4 digit octal     --
--               counter running at a frequency of 100Hz.        --
--               It is a part of the counter project. This file  --
--               contains the rtl configuration of the counter.  --
-------------------------------------------------------------------

configuration counter_rtl_cfg of counter is
	for rtl
	end for;
end counter_rtl_cfg;
